module sra(
    //input 
	 input logic [31:0] a_i,
	 input logic [4:0] b_i,
	 //output 
	 output logic [31:0]c_i);
	 always @(*) begin
	 case(b_i)
	 0: c_i <= a_i;
	 1: c_i <= {a_i[31], a_i[31:1]};
	 2: c_i <= {{2{a_i[31]}}, a_i[31:2]};
	 3: c_i <= {{3{a_i[31]}}, a_i[31:3]};
	 4: c_i <= {{4{a_i[31]}}, a_i[31:4]};
	 5: c_i <= {{5{a_i[31]}}, a_i[31:5]};
	 6: c_i <= {{6{a_i[31]}}, a_i[31:6]};
	 7: c_i <= {{7{a_i[31]}}, a_i[31:7]};
	 8: c_i <= {{8{a_i[31]}}, a_i[31:8]};
	 9: c_i <= {{9{a_i[31]}}, a_i[31:9]};
	 10: c_i <= {{10{a_i[31]}}, a_i[31:10]};
	 11: c_i <= {{11{a_i[31]}}, a_i[31:11]};
	 12: c_i <= {{12{a_i[31]}}, a_i[31:12]};
	 13: c_i <= {{13{a_i[31]}}, a_i[31:13]};
	 14: c_i <= {{14{a_i[31]}}, a_i[31:14]};
	 15: c_i <= {{15{a_i[31]}}, a_i[31:15]};
	 16: c_i <= {{16{a_i[31]}}, a_i[31:16]};
	 17: c_i <= {{17{a_i[31]}}, a_i[31:17]};
	 18: c_i <= {{18{a_i[31]}}, a_i[31:18]};
	 19: c_i <= {{19{a_i[31]}}, a_i[31:19]};
	 20: c_i <= {{20{a_i[31]}}, a_i[31:20]};
	 21: c_i <= {{21{a_i[31]}}, a_i[31:21]};
	 22: c_i <= {{22{a_i[31]}}, a_i[31:22]};
	 23: c_i <= {{23{a_i[31]}}, a_i[31:23]};
	 24: c_i <= {{24{a_i[31]}}, a_i[31:24]};
	 25: c_i <= {{25{a_i[31]}}, a_i[31:25]};
	 26: c_i <= {{26{a_i[31]}}, a_i[31:26]};
	 27: c_i <= {{27{a_i[31]}}, a_i[31:27]};
	 28: c_i <= {{28{a_i[31]}}, a_i[31:28]};
	 29: c_i <= {{29{a_i[31]}}, a_i[31:29]};
	 30: c_i <= {{30{a_i[31]}}, a_i[31:30]};
	 31: c_i <= {32{a_i[31]}};
	 endcase
	 end
endmodule 